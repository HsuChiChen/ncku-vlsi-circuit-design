* SPICE NETLIST
***************************************

.SUBCKT L POS NEG
.ENDS
***************************************
.SUBCKT tristate_inv GND D0 Y S D1 VDD
** N=11 EP=6 IP=0 FDC=10
M0 10 D0 GND GND N_18 L=1.8e-07 W=5e-07 AD=6.375e-14 AS=2.45e-13 PD=2.55e-07 PS=1.48e-06 $X=160 $Y=-1280 $D=0
M1 Y 7 10 GND N_18 L=1.8e-07 W=5e-07 AD=1.9e-13 AS=6.375e-14 PD=7.6e-07 PS=2.55e-07 $X=595 $Y=-1280 $D=0
M2 11 S Y GND N_18 L=1.8e-07 W=5e-07 AD=1.025e-13 AS=1.9e-13 PD=4.1e-07 PS=7.6e-07 $X=1535 $Y=-1280 $D=0
M3 GND D1 11 GND N_18 L=1.8e-07 W=5e-07 AD=1.3875e-13 AS=1.025e-13 PD=5.55e-07 PS=4.1e-07 $X=2125 $Y=-1280 $D=0
M4 7 S GND GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.3875e-13 PD=1.48e-06 PS=5.55e-07 $X=2860 $Y=-1280 $D=0
M5 8 D0 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=1.275e-13 AS=4.95e-13 PD=2.55e-07 PS=1.99e-06 $X=160 $Y=1095 $D=1
M6 Y S 8 VDD P_18 L=1.8e-07 W=1e-06 AD=4.425e-13 AS=1.275e-13 PD=8.85e-07 PS=2.55e-07 $X=595 $Y=1095 $D=1
M7 9 7 Y VDD P_18 L=1.8e-07 W=1e-06 AD=1.425e-13 AS=4.425e-13 PD=2.85e-07 PS=8.85e-07 $X=1660 $Y=1095 $D=1
M8 VDD D1 9 VDD P_18 L=1.8e-07 W=1e-06 AD=2.775e-13 AS=1.425e-13 PD=5.55e-07 PS=2.85e-07 $X=2125 $Y=1095 $D=1
M9 7 S VDD VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.775e-13 PD=1.98e-06 PS=5.55e-07 $X=2860 $Y=1095 $D=1
.ENDS
***************************************
