* SPICE NETLIST
***************************************

.SUBCKT L POS NEG
.ENDS
***************************************
.SUBCKT decoder_3to8 W2 W1 W0 EN Y7 Y6 Y5 Y4 Y3 Y2 Y1 Y0 GND VDD
** N=42 EP=14 IP=0 FDC=72
M0 1 EN GND GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.475e-13 PD=1.48e-06 PS=1.49e-06 $X=-41120 $Y=-2430 $D=0
M1 3 W2 GND GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.475e-13 PD=1.48e-06 PS=1.49e-06 $X=-39655 $Y=-2405 $D=0
M2 4 W2 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=-38060 $Y=-2440 $D=0
M3 GND 1 4 GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=-37370 $Y=-2440 $D=0
M4 5 3 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=-35905 $Y=-2440 $D=0
M5 GND 1 5 GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=-35215 $Y=-2440 $D=0
M6 6 5 GND GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.475e-13 PD=1.48e-06 PS=1.49e-06 $X=-33745 $Y=-2430 $D=0
M7 8 W1 GND GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.475e-13 PD=1.48e-06 PS=1.49e-06 $X=-32280 $Y=-2430 $D=0
M8 10 W0 GND GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.475e-13 PD=1.48e-06 PS=1.49e-06 $X=-30815 $Y=-2430 $D=0
M9 GND 6 Y7 GND N_18 L=1.8e-07 W=5e-07 AD=1.35e-13 AS=2.45e-13 PD=5.4e-07 PS=1.48e-06 $X=-29315 $Y=-2430 $D=0
M10 Y7 10 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.35e-13 PD=5.1e-07 PS=5.4e-07 $X=-28595 $Y=-2430 $D=0
M11 GND 8 Y7 GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=-27905 $Y=-2430 $D=0
M12 GND 6 Y6 GND N_18 L=1.8e-07 W=5e-07 AD=1.35e-13 AS=2.45e-13 PD=5.4e-07 PS=1.48e-06 $X=-26445 $Y=-2430 $D=0
M13 Y6 W0 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.35e-13 PD=5.1e-07 PS=5.4e-07 $X=-25725 $Y=-2430 $D=0
M14 GND 8 Y6 GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=-25035 $Y=-2430 $D=0
M15 GND 6 Y5 GND N_18 L=1.8e-07 W=5e-07 AD=1.35e-13 AS=2.45e-13 PD=5.4e-07 PS=1.48e-06 $X=-23570 $Y=-2430 $D=0
M16 Y5 10 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.35e-13 PD=5.1e-07 PS=5.4e-07 $X=-22850 $Y=-2430 $D=0
M17 GND W1 Y5 GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=-22160 $Y=-2430 $D=0
M18 GND 6 Y4 GND N_18 L=1.8e-07 W=5e-07 AD=1.35e-13 AS=2.45e-13 PD=5.4e-07 PS=1.48e-06 $X=-20700 $Y=-2430 $D=0
M19 Y4 W0 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.35e-13 PD=5.1e-07 PS=5.4e-07 $X=-19980 $Y=-2430 $D=0
M20 GND W1 Y4 GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=-19290 $Y=-2430 $D=0
M21 11 4 GND GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.475e-13 PD=1.48e-06 PS=1.49e-06 $X=-17820 $Y=-2430 $D=0
M22 12 W1 GND GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.475e-13 PD=1.48e-06 PS=1.49e-06 $X=-16355 $Y=-2430 $D=0
M23 13 W0 GND GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.475e-13 PD=1.48e-06 PS=1.49e-06 $X=-14890 $Y=-2430 $D=0
M24 GND 11 Y3 GND N_18 L=1.8e-07 W=5e-07 AD=1.35e-13 AS=2.45e-13 PD=5.4e-07 PS=1.48e-06 $X=-13390 $Y=-2430 $D=0
M25 Y3 13 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.35e-13 PD=5.1e-07 PS=5.4e-07 $X=-12670 $Y=-2430 $D=0
M26 GND 12 Y3 GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=-11980 $Y=-2430 $D=0
M27 GND 11 Y2 GND N_18 L=1.8e-07 W=5e-07 AD=1.35e-13 AS=2.45e-13 PD=5.4e-07 PS=1.48e-06 $X=-10520 $Y=-2430 $D=0
M28 Y2 W0 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.35e-13 PD=5.1e-07 PS=5.4e-07 $X=-9800 $Y=-2430 $D=0
M29 GND 12 Y2 GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=-9110 $Y=-2430 $D=0
M30 GND 11 Y1 GND N_18 L=1.8e-07 W=5e-07 AD=1.35e-13 AS=2.45e-13 PD=5.4e-07 PS=1.48e-06 $X=-7645 $Y=-2430 $D=0
M31 Y1 13 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.35e-13 PD=5.1e-07 PS=5.4e-07 $X=-6925 $Y=-2430 $D=0
M32 GND W1 Y1 GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=-6235 $Y=-2430 $D=0
M33 GND 11 Y0 GND N_18 L=1.8e-07 W=5e-07 AD=1.35e-13 AS=2.45e-13 PD=5.4e-07 PS=1.48e-06 $X=-4775 $Y=-2430 $D=0
M34 Y0 W0 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.35e-13 PD=5.1e-07 PS=5.4e-07 $X=-4055 $Y=-2430 $D=0
M35 GND W1 Y0 GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=-3365 $Y=-2430 $D=0
M36 1 EN VDD VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06 $X=-41120 $Y=-795 $D=1
M37 3 W2 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06 $X=-39655 $Y=-770 $D=1
M38 25 W2 4 VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06 $X=-38060 $Y=-805 $D=1
M39 VDD 1 25 VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07 $X=-37370 $Y=-805 $D=1
M40 26 3 5 VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06 $X=-35905 $Y=-805 $D=1
M41 VDD 1 26 VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07 $X=-35215 $Y=-805 $D=1
M42 6 5 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06 $X=-33745 $Y=-795 $D=1
M43 8 W1 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06 $X=-32280 $Y=-795 $D=1
M44 10 W0 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06 $X=-30815 $Y=-795 $D=1
M45 27 6 Y7 VDD P_18 L=1.8e-07 W=1e-06 AD=2.7e-13 AS=4.9e-13 PD=5.4e-07 PS=1.98e-06 $X=-29315 $Y=-795 $D=1
M46 28 10 27 VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=2.7e-13 PD=5.1e-07 PS=5.4e-07 $X=-28595 $Y=-795 $D=1
M47 VDD 8 28 VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07 $X=-27905 $Y=-795 $D=1
M48 29 6 Y6 VDD P_18 L=1.8e-07 W=1e-06 AD=2.7e-13 AS=4.9e-13 PD=5.4e-07 PS=1.98e-06 $X=-26445 $Y=-795 $D=1
M49 30 W0 29 VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=2.7e-13 PD=5.1e-07 PS=5.4e-07 $X=-25725 $Y=-795 $D=1
M50 VDD 8 30 VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07 $X=-25035 $Y=-795 $D=1
M51 31 6 Y5 VDD P_18 L=1.8e-07 W=1e-06 AD=2.7e-13 AS=4.9e-13 PD=5.4e-07 PS=1.98e-06 $X=-23570 $Y=-795 $D=1
M52 32 10 31 VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=2.7e-13 PD=5.1e-07 PS=5.4e-07 $X=-22850 $Y=-795 $D=1
M53 VDD W1 32 VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07 $X=-22160 $Y=-795 $D=1
M54 33 6 Y4 VDD P_18 L=1.8e-07 W=1e-06 AD=2.7e-13 AS=4.9e-13 PD=5.4e-07 PS=1.98e-06 $X=-20700 $Y=-795 $D=1
M55 34 W0 33 VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=2.7e-13 PD=5.1e-07 PS=5.4e-07 $X=-19980 $Y=-795 $D=1
M56 VDD W1 34 VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07 $X=-19290 $Y=-795 $D=1
M57 11 4 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06 $X=-17820 $Y=-795 $D=1
M58 12 W1 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06 $X=-16355 $Y=-795 $D=1
M59 13 W0 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06 $X=-14890 $Y=-795 $D=1
M60 35 11 Y3 VDD P_18 L=1.8e-07 W=1e-06 AD=2.7e-13 AS=4.9e-13 PD=5.4e-07 PS=1.98e-06 $X=-13390 $Y=-795 $D=1
M61 36 13 35 VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=2.7e-13 PD=5.1e-07 PS=5.4e-07 $X=-12670 $Y=-795 $D=1
M62 VDD 12 36 VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07 $X=-11980 $Y=-795 $D=1
M63 37 11 Y2 VDD P_18 L=1.8e-07 W=1e-06 AD=2.7e-13 AS=4.9e-13 PD=5.4e-07 PS=1.98e-06 $X=-10520 $Y=-795 $D=1
M64 38 W0 37 VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=2.7e-13 PD=5.1e-07 PS=5.4e-07 $X=-9800 $Y=-795 $D=1
M65 VDD 12 38 VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07 $X=-9110 $Y=-795 $D=1
M66 39 11 Y1 VDD P_18 L=1.8e-07 W=1e-06 AD=2.7e-13 AS=4.9e-13 PD=5.4e-07 PS=1.98e-06 $X=-7645 $Y=-795 $D=1
M67 40 13 39 VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=2.7e-13 PD=5.1e-07 PS=5.4e-07 $X=-6925 $Y=-795 $D=1
M68 VDD W1 40 VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07 $X=-6235 $Y=-795 $D=1
M69 41 11 Y0 VDD P_18 L=1.8e-07 W=1e-06 AD=2.7e-13 AS=4.9e-13 PD=5.4e-07 PS=1.98e-06 $X=-4775 $Y=-795 $D=1
M70 42 W0 41 VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=2.7e-13 PD=5.1e-07 PS=5.4e-07 $X=-4055 $Y=-795 $D=1
M71 VDD W1 42 VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07 $X=-3365 $Y=-795 $D=1
.ENDS
***************************************
