************************************************************************
* auCdl Netlist:
* 
* Library Name:  lab
* Top Cell Name: inv
* View Name:     schematic
* Netlisted on:  Mar 31 16:31:22 2022
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: lab
* Cell Name:    inv
* View Name:    schematic
************************************************************************

.SUBCKT inv GND VDD in out
*.PININFO GND:I VDD:I in:I out:O
MM5 out in GND GND n_18 W=2u L=180.00n
MM4 out in VDD VDD p_18 W=6u L=180.00n
.ENDS

