* SPICE NETLIST
***************************************

.SUBCKT L POS NEG
.ENDS
***************************************
.SUBCKT aoi31 D A Y B C GND VDD
** N=10 EP=7 IP=0 FDC=8
M0 Y D GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=-380 $Y=-2210 $D=0
M1 9 A Y GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=310 $Y=-2210 $D=0
M2 10 B 9 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=1000 $Y=-2210 $D=0
M3 GND C 10 GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=1690 $Y=-2210 $D=0
M4 5 D Y VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06 $X=-380 $Y=-505 $D=1
M5 VDD A 5 VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=2.55e-13 PD=5.1e-07 PS=5.1e-07 $X=310 $Y=-505 $D=1
M6 5 B VDD VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=2.55e-13 PD=5.1e-07 PS=5.1e-07 $X=1000 $Y=-505 $D=1
M7 VDD C 5 VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07 $X=1690 $Y=-505 $D=1
.ENDS
***************************************
