* SPICE NETLIST
***************************************

.SUBCKT L POS NEG
.ENDS
***************************************
.SUBCKT ring_oscillator vin GND VDD
** N=7 EP=3 IP=0 FDC=20
M0 1 vin GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=1505 $Y=-1005 $D=0
M1 GND vin 1 GND N_18 L=1.8e-07 W=5e-07 AD=1.425e-13 AS=1.275e-13 PD=5.7e-07 PS=5.1e-07 $X=2195 $Y=-1005 $D=0
M2 2 1 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.425e-13 PD=5.1e-07 PS=5.7e-07 $X=2945 $Y=-1005 $D=0
M3 GND 1 2 GND N_18 L=1.8e-07 W=5e-07 AD=1.425e-13 AS=1.275e-13 PD=5.7e-07 PS=5.1e-07 $X=3635 $Y=-1005 $D=0
M4 3 2 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.425e-13 PD=5.1e-07 PS=5.7e-07 $X=4385 $Y=-1005 $D=0
M5 GND 2 3 GND N_18 L=1.8e-07 W=5e-07 AD=1.425e-13 AS=1.275e-13 PD=5.7e-07 PS=5.1e-07 $X=5075 $Y=-1005 $D=0
M6 4 3 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.425e-13 PD=5.1e-07 PS=5.7e-07 $X=5825 $Y=-1005 $D=0
M7 GND 3 4 GND N_18 L=1.8e-07 W=5e-07 AD=1.425e-13 AS=1.275e-13 PD=5.7e-07 PS=5.1e-07 $X=6515 $Y=-1005 $D=0
M8 vin 4 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.425e-13 PD=5.1e-07 PS=5.7e-07 $X=7265 $Y=-1005 $D=0
M9 GND 4 vin GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=7955 $Y=-1005 $D=0
M10 1 vin VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13 AS=7.35e-13 PD=5.1e-07 PS=2.48e-06 $X=1505 $Y=475 $D=1
M11 VDD vin 1 VDD P_18 L=1.8e-07 W=1.5e-06 AD=4.275e-13 AS=3.825e-13 PD=5.7e-07 PS=5.1e-07 $X=2195 $Y=475 $D=1
M12 2 1 VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13 AS=4.275e-13 PD=5.1e-07 PS=5.7e-07 $X=2945 $Y=475 $D=1
M13 VDD 1 2 VDD P_18 L=1.8e-07 W=1.5e-06 AD=4.275e-13 AS=3.825e-13 PD=5.7e-07 PS=5.1e-07 $X=3635 $Y=475 $D=1
M14 3 2 VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13 AS=4.275e-13 PD=5.1e-07 PS=5.7e-07 $X=4385 $Y=475 $D=1
M15 VDD 2 3 VDD P_18 L=1.8e-07 W=1.5e-06 AD=4.275e-13 AS=3.825e-13 PD=5.7e-07 PS=5.1e-07 $X=5075 $Y=475 $D=1
M16 4 3 VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13 AS=4.275e-13 PD=5.1e-07 PS=5.7e-07 $X=5825 $Y=475 $D=1
M17 VDD 3 4 VDD P_18 L=1.8e-07 W=1.5e-06 AD=4.275e-13 AS=3.825e-13 PD=5.7e-07 PS=5.1e-07 $X=6515 $Y=475 $D=1
M18 vin 4 VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13 AS=4.275e-13 PD=5.1e-07 PS=5.7e-07 $X=7265 $Y=475 $D=1
M19 VDD 4 vin VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=3.825e-13 PD=2.48e-06 PS=5.1e-07 $X=7955 $Y=475 $D=1
.ENDS
***************************************
