************************************************************************
* auCdl Netlist:
* 
* Library Name:  lab1
* Top Cell Name: decoder_3to8
* View Name:     schematic
* Netlisted on:  Mar 25 21:07:21 2022
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: lab1
* Cell Name:    nor
* View Name:    schematic
************************************************************************

.SUBCKT nor A B GND VDD Y
*.PININFO A:I B:I GND:I VDD:I Y:O
MM1 Y B net4 VDD p_18 W=1u L=180.00n
MM0 net4 A VDD VDD p_18 W=1u L=180.00n
MM6 Y B GND GND n_18 W=500.0n L=180.00n
MM5 Y A GND GND n_18 W=500.0n L=180.00n
.ENDS

************************************************************************
* Library Name: lab1
* Cell Name:    inv
* View Name:    schematic
************************************************************************

.SUBCKT inv GND VDD in out
*.PININFO GND:I VDD:I in:I out:O
MM5 out in GND GND n_18 W=500.0n L=180.00n
MM4 out in VDD VDD p_18 W=1u L=180.00n
.ENDS

************************************************************************
* Library Name: lab1
* Cell Name:    nor_3
* View Name:    schematic
************************************************************************

.SUBCKT nor_3 A B C GND VDD Y
*.PININFO A:I B:I C:I GND:I VDD:I Y:O
MM2 Y C net1 VDD p_18 W=1u L=180.00n
MM1 net1 B net4 VDD p_18 W=1u L=180.00n
MM0 net4 A VDD VDD p_18 W=1u L=180.00n
MM8 Y C GND GND n_18 W=500.0n L=180.00n
MM6 Y B GND GND n_18 W=500.0n L=180.00n
MM5 Y A GND GND n_18 W=500.0n L=180.00n
.ENDS

************************************************************************
* Library Name: lab1
* Cell Name:    decoder_2to4
* View Name:    schematic
************************************************************************

.SUBCKT decoder_2to4 EN GND VDD W0 W1 Y0 Y1 Y2 Y3
*.PININFO EN:I GND:I VDD:I W0:I W1:I Y0:O Y1:O Y2:O Y3:O
XI7 GND VDD EN net1 / inv
XI1 GND VDD W0 net6 / inv
XI0 GND VDD W1 net4 / inv
XI2 W0 net1 W1 GND VDD Y0 / nor_3
XI3 net6 net1 W1 GND VDD Y1 / nor_3
XI4 W0 net1 net4 GND VDD Y2 / nor_3
XI5 net6 net1 net4 GND VDD Y3 / nor_3
.ENDS

************************************************************************
* Library Name: lab1
* Cell Name:    decoder_3to8
* View Name:    schematic
************************************************************************

.SUBCKT decoder_3to8 EN GND VDD W0 W1 W2 Y0 Y1 Y2 Y3 Y4 Y5 Y6 Y7
*.PININFO EN:I GND:I VDD:I W0:I W1:I W2:I Y0:O Y1:O Y2:O Y3:O Y4:O Y5:O Y6:O 
*.PININFO Y7:O
XI3 net19 net15 GND VDD net6 / nor
XI2 W2 net15 GND VDD net1 / nor
XI5 GND VDD EN net15 / inv
XI4 GND VDD W2 net19 / inv
XI1 net6 GND VDD W0 W1 Y4 Y5 Y6 Y7 / decoder_2to4
XI0 net1 GND VDD W0 W1 Y0 Y1 Y2 Y3 / decoder_2to4
.ENDS

