************************************************************************
* auCdl Netlist:
* 
* Library Name:  lab
* Top Cell Name: path_delay_1
* View Name:     schematic
* Netlisted on:  Apr  8 21:27:30 2022
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: lab
* Cell Name:    nand_6
* View Name:    schematic
************************************************************************

.SUBCKT nand_6 A B C D E F GND VDD Y
*.PININFO A:I B:I C:I D:I E:I F:I GND:I VDD:I Y:O
MM13 Y F VDD VDD p_18 W=1.25u L=180.00n
MM8 Y E VDD VDD p_18 W=1.25u L=180.00n
MM7 Y D VDD VDD p_18 W=1.25u L=180.00n
MM4 Y C VDD VDD p_18 W=1.25u L=180.00n
MM1 Y B VDD VDD p_18 W=1.25u L=180.00n
MM0 Y A VDD VDD p_18 W=1.25u L=180.00n
MM12 net11 F GND GND n_18 W=3.75u L=180.00n
MM11 net3 E net11 GND n_18 W=3.75u L=180.00n
MM10 net2 D net3 GND n_18 W=3.75u L=180.00n
MM6 net1 B net4 GND n_18 W=3.75u L=180.00n
MM5 Y A net1 GND n_18 W=3.75u L=180.00n
MM9 net4 C net2 GND n_18 W=3.75u L=180.00n
.ENDS

************************************************************************
* Library Name: lab
* Cell Name:    inv
* View Name:    schematic
************************************************************************

.SUBCKT inv GND VDD in out
*.PININFO GND:I VDD:I in:I out:O
MM5 out in GND GND n_18 W=10.21u L=180.00n
MM4 out in VDD VDD p_18 W=20.42u L=180.00n
.ENDS

************************************************************************
* Library Name: lab
* Cell Name:    path_delay_1
* View Name:    schematic
************************************************************************

.SUBCKT path_delay_1 GND VDD out pulse_in
*.PININFO GND:I VDD:I pulse_in:I out:O
XI0 VDD VDD VDD VDD VDD pulse_in GND VDD net1 / nand_6
XI8 GND VDD net1 out / inv
.ENDS

