* SPICE NETLIST
***************************************

.SUBCKT L POS NEG
.ENDS
***************************************
.SUBCKT d_latch Q CLK D VDD GND Q_INV
** N=8 EP=6 IP=0 FDC=10
M0 6 7 Q GND N_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06 $X=-1290 $Y=-3925 $D=0
M1 D CLK Q GND N_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06 $X=-1290 $Y=1280 $D=0
M2 7 CLK GND GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=1915 $Y=1720 $D=0
M3 GND Q_INV 6 GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=2560 $Y=-7395 $D=0
M4 GND Q Q_INV GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=4565 $Y=-7395 $D=0
M5 6 CLK Q VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06 $X=-1290 $Y=-6065 $D=1
M6 D 7 Q VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06 $X=-1290 $Y=-860 $D=1
M7 7 CLK VDD VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06 $X=1915 $Y=3825 $D=1
M8 VDD Q_INV 6 VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06 $X=2560 $Y=-5290 $D=1
M9 VDD Q Q_INV VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06 $X=4565 $Y=-5290 $D=1
.ENDS
***************************************
