* SPICE NETLIST
***************************************

.SUBCKT L POS NEG
.ENDS
***************************************
.SUBCKT path_delay_4 out GND pulse_in VDD
** N=14 EP=4 IP=0 FDC=60
M0 3 1 4 GND N_18 L=1.8e-07 W=4.47e-06 AD=1.13985e-12 AS=2.1903e-12 PD=5.1e-07 PS=5.45e-06 $X=-18715 $Y=-7220 $D=0
M1 4 1 3 GND N_18 L=1.8e-07 W=4.47e-06 AD=1.13985e-12 AS=1.13985e-12 PD=5.1e-07 PS=5.1e-07 $X=-18025 $Y=-7220 $D=0
M2 3 1 4 GND N_18 L=1.8e-07 W=4.47e-06 AD=1.13985e-12 AS=1.13985e-12 PD=5.1e-07 PS=5.1e-07 $X=-17335 $Y=-7220 $D=0
M3 4 1 3 GND N_18 L=1.8e-07 W=4.47e-06 AD=1.13985e-12 AS=1.13985e-12 PD=5.1e-07 PS=5.1e-07 $X=-16645 $Y=-7220 $D=0
M4 3 1 4 GND N_18 L=1.8e-07 W=4.47e-06 AD=1.13985e-12 AS=1.13985e-12 PD=5.1e-07 PS=5.1e-07 $X=-15955 $Y=-7220 $D=0
M5 GND 2 3 GND N_18 L=1.8e-07 W=4.47e-06 AD=1.13985e-12 AS=1.13985e-12 PD=5.1e-07 PS=5.1e-07 $X=-15265 $Y=-7220 $D=0
M6 3 2 GND GND N_18 L=1.8e-07 W=4.47e-06 AD=1.13985e-12 AS=1.13985e-12 PD=5.1e-07 PS=5.1e-07 $X=-14575 $Y=-7220 $D=0
M7 GND 2 3 GND N_18 L=1.8e-07 W=4.47e-06 AD=1.13985e-12 AS=1.13985e-12 PD=5.1e-07 PS=5.1e-07 $X=-13885 $Y=-7220 $D=0
M8 3 2 GND GND N_18 L=1.8e-07 W=4.47e-06 AD=1.13985e-12 AS=1.13985e-12 PD=5.1e-07 PS=5.1e-07 $X=-13195 $Y=-7220 $D=0
M9 GND 2 3 GND N_18 L=1.8e-07 W=4.47e-06 AD=1.13265e-12 AS=1.13985e-12 PD=7.88225e-07 PS=5.1e-07 $X=-12505 $Y=-7220 $D=0
M10 out 4 GND GND N_18 L=1.8e-07 W=4.32e-06 AD=1.1016e-12 AS=1.09465e-12 PD=5.1e-07 PS=7.61775e-07 $X=-11815 $Y=-6880 $D=0
M11 GND 4 out GND N_18 L=1.8e-07 W=4.32e-06 AD=1.1016e-12 AS=1.1016e-12 PD=5.1e-07 PS=5.1e-07 $X=-11125 $Y=-6880 $D=0
M12 out 4 GND GND N_18 L=1.8e-07 W=4.32e-06 AD=1.1016e-12 AS=1.1016e-12 PD=5.1e-07 PS=5.1e-07 $X=-10435 $Y=-6880 $D=0
M13 GND 4 out GND N_18 L=1.8e-07 W=4.32e-06 AD=1.1016e-12 AS=1.1016e-12 PD=5.1e-07 PS=5.1e-07 $X=-9745 $Y=-6880 $D=0
M14 out 4 GND GND N_18 L=1.8e-07 W=4.32e-06 AD=1.1016e-12 AS=1.1016e-12 PD=5.1e-07 PS=5.1e-07 $X=-9055 $Y=-6880 $D=0
M15 GND 4 out GND N_18 L=1.8e-07 W=4.32e-06 AD=1.1016e-12 AS=1.1016e-12 PD=5.1e-07 PS=5.1e-07 $X=-8365 $Y=-6880 $D=0
M16 out 4 GND GND N_18 L=1.8e-07 W=4.32e-06 AD=1.1016e-12 AS=1.1016e-12 PD=5.1e-07 PS=5.1e-07 $X=-7675 $Y=-6880 $D=0
M17 GND 4 out GND N_18 L=1.8e-07 W=4.32e-06 AD=1.1016e-12 AS=1.1016e-12 PD=5.1e-07 PS=5.1e-07 $X=-6985 $Y=-6880 $D=0
M18 out 4 GND GND N_18 L=1.8e-07 W=4.32e-06 AD=1.1016e-12 AS=1.1016e-12 PD=5.1e-07 PS=5.1e-07 $X=-6295 $Y=-6880 $D=0
M19 GND 4 out GND N_18 L=1.8e-07 W=4.32e-06 AD=2.1168e-12 AS=1.1016e-12 PD=5.3e-06 PS=5.1e-07 $X=-5605 $Y=-6880 $D=0
M20 11 VDD 6 GND N_18 L=1.8e-07 W=3e-06 AD=3.75e-13 AS=1.47e-12 PD=2.5e-07 PS=3.98e-06 $X=-2180 $Y=-1475 $D=0
M21 12 VDD 11 GND N_18 L=1.8e-07 W=3e-06 AD=3.75e-13 AS=3.75e-13 PD=2.5e-07 PS=2.5e-07 $X=-1750 $Y=-1475 $D=0
M22 GND VDD 12 GND N_18 L=1.8e-07 W=3e-06 AD=6.44544e-13 AS=3.75e-13 PD=1.27181e-06 PS=2.5e-07 $X=-1320 $Y=-1475 $D=0
M23 1 6 GND GND N_18 L=1.8e-07 W=1.93e-06 AD=4.9215e-13 AS=4.14656e-13 PD=5.1e-07 PS=8.18195e-07 $X=-630 $Y=-405 $D=0
M24 GND 6 1 GND N_18 L=1.8e-07 W=1.93e-06 AD=4.9215e-13 AS=4.9215e-13 PD=5.1e-07 PS=5.1e-07 $X=60 $Y=-405 $D=0
M25 2 9 GND GND N_18 L=1.8e-07 W=1.93e-06 AD=4.9215e-13 AS=4.9215e-13 PD=5.1e-07 PS=5.1e-07 $X=750 $Y=-405 $D=0
M26 GND 9 2 GND N_18 L=1.8e-07 W=1.93e-06 AD=4.14656e-13 AS=4.9215e-13 PD=8.18195e-07 PS=5.1e-07 $X=1440 $Y=-405 $D=0
M27 13 pulse_in GND GND N_18 L=1.8e-07 W=3e-06 AD=3.75e-13 AS=6.44544e-13 PD=2.5e-07 PS=1.27181e-06 $X=2130 $Y=-1475 $D=0
M28 14 VDD 13 GND N_18 L=1.8e-07 W=3e-06 AD=3.75e-13 AS=3.75e-13 PD=2.5e-07 PS=2.5e-07 $X=2560 $Y=-1475 $D=0
M29 9 VDD 14 GND N_18 L=1.8e-07 W=3e-06 AD=1.47e-12 AS=3.75e-13 PD=3.98e-06 PS=2.5e-07 $X=2990 $Y=-1475 $D=0
M30 VDD 1 4 VDD P_18 L=1.8e-07 W=7.45e-06 AD=1.89975e-12 AS=3.6505e-12 PD=5.1e-07 PS=8.43e-06 $X=-17335 $Y=-1630 $D=1
M31 4 1 VDD VDD P_18 L=1.8e-07 W=7.45e-06 AD=1.89975e-12 AS=1.89975e-12 PD=5.1e-07 PS=5.1e-07 $X=-16645 $Y=-1630 $D=1
M32 VDD 1 4 VDD P_18 L=1.8e-07 W=7.45e-06 AD=1.89975e-12 AS=1.89975e-12 PD=5.1e-07 PS=5.1e-07 $X=-15955 $Y=-1630 $D=1
M33 4 2 VDD VDD P_18 L=1.8e-07 W=7.45e-06 AD=1.89975e-12 AS=1.89975e-12 PD=5.1e-07 PS=5.1e-07 $X=-15265 $Y=-1630 $D=1
M34 VDD 2 4 VDD P_18 L=1.8e-07 W=7.45e-06 AD=1.89975e-12 AS=1.89975e-12 PD=5.1e-07 PS=5.1e-07 $X=-14575 $Y=-1630 $D=1
M35 4 2 VDD VDD P_18 L=1.8e-07 W=7.45e-06 AD=3.6505e-12 AS=1.89975e-12 PD=8.43e-06 PS=5.1e-07 $X=-13885 $Y=-1630 $D=1
M36 out 4 VDD VDD P_18 L=1.8e-07 W=8.64e-06 AD=2.2032e-12 AS=4.2336e-12 PD=5.1e-07 PS=9.62e-06 $X=-11815 $Y=-1630 $D=1
M37 VDD 4 out VDD P_18 L=1.8e-07 W=8.64e-06 AD=2.2032e-12 AS=2.2032e-12 PD=5.1e-07 PS=5.1e-07 $X=-11125 $Y=-1630 $D=1
M38 out 4 VDD VDD P_18 L=1.8e-07 W=8.64e-06 AD=2.2032e-12 AS=2.2032e-12 PD=5.1e-07 PS=5.1e-07 $X=-10435 $Y=-1630 $D=1
M39 VDD 4 out VDD P_18 L=1.8e-07 W=8.64e-06 AD=2.2032e-12 AS=2.2032e-12 PD=5.1e-07 PS=5.1e-07 $X=-9745 $Y=-1630 $D=1
M40 out 4 VDD VDD P_18 L=1.8e-07 W=8.64e-06 AD=2.2032e-12 AS=2.2032e-12 PD=5.1e-07 PS=5.1e-07 $X=-9055 $Y=-1630 $D=1
M41 VDD 4 out VDD P_18 L=1.8e-07 W=8.64e-06 AD=2.2032e-12 AS=2.2032e-12 PD=5.1e-07 PS=5.1e-07 $X=-8365 $Y=-1630 $D=1
M42 out 4 VDD VDD P_18 L=1.8e-07 W=8.64e-06 AD=2.2032e-12 AS=2.2032e-12 PD=5.1e-07 PS=5.1e-07 $X=-7675 $Y=-1630 $D=1
M43 VDD 4 out VDD P_18 L=1.8e-07 W=8.64e-06 AD=2.2032e-12 AS=2.2032e-12 PD=5.1e-07 PS=5.1e-07 $X=-6985 $Y=-1630 $D=1
M44 out 4 VDD VDD P_18 L=1.8e-07 W=8.64e-06 AD=2.2032e-12 AS=2.2032e-12 PD=5.1e-07 PS=5.1e-07 $X=-6295 $Y=-1630 $D=1
M45 VDD 4 out VDD P_18 L=1.8e-07 W=8.64e-06 AD=4.2336e-12 AS=2.2032e-12 PD=9.62e-06 PS=5.1e-07 $X=-5605 $Y=-1630 $D=1
M46 VDD VDD 6 VDD P_18 L=1.8e-07 W=2e-06 AD=5.1e-13 AS=9.8e-13 PD=5.1e-07 PS=2.98e-06 $X=-4145 $Y=3980 $D=1
M47 6 VDD VDD VDD P_18 L=1.8e-07 W=2e-06 AD=5.1e-13 AS=5.1e-13 PD=5.1e-07 PS=5.1e-07 $X=-3455 $Y=3980 $D=1
M48 VDD VDD 6 VDD P_18 L=1.8e-07 W=2e-06 AD=5.11603e-13 AS=5.1e-13 PD=5.54707e-07 PS=5.1e-07 $X=-2765 $Y=3980 $D=1
M49 1 6 VDD VDD P_18 L=1.8e-07 W=1.93e-06 AD=5.54875e-13 AS=4.93697e-13 PD=5.75e-07 PS=5.35293e-07 $X=-2075 $Y=3980 $D=1
M50 VDD 6 1 VDD P_18 L=1.8e-07 W=1.93e-06 AD=4.9215e-13 AS=5.54875e-13 PD=5.1e-07 PS=5.75e-07 $X=-1320 $Y=3980 $D=1
M51 1 6 VDD VDD P_18 L=1.8e-07 W=1.93e-06 AD=4.9215e-13 AS=4.9215e-13 PD=5.1e-07 PS=5.1e-07 $X=-630 $Y=3980 $D=1
M52 VDD 6 1 VDD P_18 L=1.8e-07 W=1.93e-06 AD=4.9215e-13 AS=4.9215e-13 PD=5.1e-07 PS=5.1e-07 $X=60 $Y=3980 $D=1
M53 2 9 VDD VDD P_18 L=1.8e-07 W=1.93e-06 AD=4.9215e-13 AS=4.9215e-13 PD=5.1e-07 PS=5.1e-07 $X=750 $Y=3980 $D=1
M54 VDD 9 2 VDD P_18 L=1.8e-07 W=1.93e-06 AD=4.9215e-13 AS=4.9215e-13 PD=5.1e-07 PS=5.1e-07 $X=1440 $Y=3980 $D=1
M55 2 9 VDD VDD P_18 L=1.8e-07 W=1.93e-06 AD=5.54875e-13 AS=4.9215e-13 PD=5.75e-07 PS=5.1e-07 $X=2130 $Y=3980 $D=1
M56 VDD 9 2 VDD P_18 L=1.8e-07 W=1.93e-06 AD=4.93697e-13 AS=5.54875e-13 PD=5.35293e-07 PS=5.75e-07 $X=2885 $Y=3980 $D=1
M57 9 pulse_in VDD VDD P_18 L=1.8e-07 W=2e-06 AD=5.1e-13 AS=5.11603e-13 PD=5.1e-07 PS=5.54707e-07 $X=3575 $Y=3980 $D=1
M58 VDD VDD 9 VDD P_18 L=1.8e-07 W=2e-06 AD=5.1e-13 AS=5.1e-13 PD=5.1e-07 PS=5.1e-07 $X=4265 $Y=3980 $D=1
M59 9 VDD VDD VDD P_18 L=1.8e-07 W=2e-06 AD=9.8e-13 AS=5.1e-13 PD=2.98e-06 PS=5.1e-07 $X=4955 $Y=3980 $D=1
.ENDS
***************************************
