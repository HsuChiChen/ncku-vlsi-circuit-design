* SPICE NETLIST
***************************************

.SUBCKT L POS NEG
.ENDS
***************************************
.SUBCKT decoder_2to4 W1 W0 EN Y3 Y2 Y1 Y0 GND VDD
** N=20 EP=9 IP=0 FDC=30
M0 1 EN GND GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.475e-13 PD=1.48e-06 PS=1.49e-06 $X=-17820 $Y=-2430 $D=0
M1 3 W1 GND GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.475e-13 PD=1.48e-06 PS=1.49e-06 $X=-16355 $Y=-2430 $D=0
M2 5 W0 GND GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.475e-13 PD=1.48e-06 PS=1.49e-06 $X=-14890 $Y=-2430 $D=0
M3 GND 1 Y3 GND N_18 L=1.8e-07 W=5e-07 AD=1.35e-13 AS=2.45e-13 PD=5.4e-07 PS=1.48e-06 $X=-13390 $Y=-2430 $D=0
M4 Y3 5 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.35e-13 PD=5.1e-07 PS=5.4e-07 $X=-12670 $Y=-2430 $D=0
M5 GND 3 Y3 GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=-11980 $Y=-2430 $D=0
M6 GND 1 Y2 GND N_18 L=1.8e-07 W=5e-07 AD=1.35e-13 AS=2.45e-13 PD=5.4e-07 PS=1.48e-06 $X=-10520 $Y=-2430 $D=0
M7 Y2 W0 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.35e-13 PD=5.1e-07 PS=5.4e-07 $X=-9800 $Y=-2430 $D=0
M8 GND 3 Y2 GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=-9110 $Y=-2430 $D=0
M9 GND 1 Y1 GND N_18 L=1.8e-07 W=5e-07 AD=1.35e-13 AS=2.45e-13 PD=5.4e-07 PS=1.48e-06 $X=-7645 $Y=-2430 $D=0
M10 Y1 5 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.35e-13 PD=5.1e-07 PS=5.4e-07 $X=-6925 $Y=-2430 $D=0
M11 GND W1 Y1 GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=-6235 $Y=-2430 $D=0
M12 GND 1 Y0 GND N_18 L=1.8e-07 W=5e-07 AD=1.35e-13 AS=2.45e-13 PD=5.4e-07 PS=1.48e-06 $X=-4775 $Y=-2430 $D=0
M13 Y0 W0 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.35e-13 PD=5.1e-07 PS=5.4e-07 $X=-4055 $Y=-2430 $D=0
M14 GND W1 Y0 GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=-3365 $Y=-2430 $D=0
M15 1 EN VDD VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06 $X=-17820 $Y=-795 $D=1
M16 3 W1 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06 $X=-16355 $Y=-795 $D=1
M17 5 W0 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06 $X=-14890 $Y=-795 $D=1
M18 13 1 Y3 VDD P_18 L=1.8e-07 W=1e-06 AD=2.7e-13 AS=4.9e-13 PD=5.4e-07 PS=1.98e-06 $X=-13390 $Y=-795 $D=1
M19 14 5 13 VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=2.7e-13 PD=5.1e-07 PS=5.4e-07 $X=-12670 $Y=-795 $D=1
M20 VDD 3 14 VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07 $X=-11980 $Y=-795 $D=1
M21 15 1 Y2 VDD P_18 L=1.8e-07 W=1e-06 AD=2.7e-13 AS=4.9e-13 PD=5.4e-07 PS=1.98e-06 $X=-10520 $Y=-795 $D=1
M22 16 W0 15 VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=2.7e-13 PD=5.1e-07 PS=5.4e-07 $X=-9800 $Y=-795 $D=1
M23 VDD 3 16 VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07 $X=-9110 $Y=-795 $D=1
M24 17 1 Y1 VDD P_18 L=1.8e-07 W=1e-06 AD=2.7e-13 AS=4.9e-13 PD=5.4e-07 PS=1.98e-06 $X=-7645 $Y=-795 $D=1
M25 18 5 17 VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=2.7e-13 PD=5.1e-07 PS=5.4e-07 $X=-6925 $Y=-795 $D=1
M26 VDD W1 18 VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07 $X=-6235 $Y=-795 $D=1
M27 19 1 Y0 VDD P_18 L=1.8e-07 W=1e-06 AD=2.7e-13 AS=4.9e-13 PD=5.4e-07 PS=1.98e-06 $X=-4775 $Y=-795 $D=1
M28 20 W0 19 VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=2.7e-13 PD=5.1e-07 PS=5.4e-07 $X=-4055 $Y=-795 $D=1
M29 VDD W1 20 VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07 $X=-3365 $Y=-795 $D=1
.ENDS
***************************************
