* SPICE NETLIST
***************************************

.SUBCKT L POS NEG
.ENDS
***************************************
.SUBCKT oai14 A Y B C D VDD GND E
** N=12 EP=8 IP=0 FDC=10
M0 9 A Y GND N_18 L=1.8e-07 W=1e-06 AD=3.15e-13 AS=4.9e-13 PD=6.3e-07 PS=1.98e-06 $X=-1190 $Y=-3215 $D=0
M1 GND B 9 GND N_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=3.15e-13 PD=5.1e-07 PS=6.3e-07 $X=-380 $Y=-3215 $D=0
M2 9 C GND GND N_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=2.55e-13 PD=5.1e-07 PS=5.1e-07 $X=310 $Y=-3215 $D=0
M3 GND D 9 GND N_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=2.55e-13 PD=5.1e-07 PS=5.1e-07 $X=1000 $Y=-3215 $D=0
M4 9 E GND GND N_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07 $X=1690 $Y=-3215 $D=0
M5 Y A VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=2.46177e-13 AS=7.3255e-13 PD=1.15015e-06 PS=2.475e-06 $X=-1190 $Y=-450 $D=1
M6 10 B Y VDD P_18 L=1.8e-07 W=6e-06 AD=7.50625e-13 AS=9.88823e-13 PD=2.5e-07 PS=4.61985e-06 $X=-380 $Y=-450 $D=1
M7 11 C 10 VDD P_18 L=1.8e-07 W=6e-06 AD=7.50625e-13 AS=7.50625e-13 PD=2.5e-07 PS=2.5e-07 $X=50 $Y=-450 $D=1
M8 12 D 11 VDD P_18 L=1.8e-07 W=6e-06 AD=7.50625e-13 AS=7.50625e-13 PD=2.5e-07 PS=2.5e-07 $X=480 $Y=-450 $D=1
M9 VDD E 12 VDD P_18 L=1.8e-07 W=6e-06 AD=2.94245e-12 AS=7.50625e-13 PD=6.985e-06 PS=2.5e-07 $X=910 $Y=-450 $D=1
.ENDS
***************************************
