* SPICE NETLIST
***************************************

.SUBCKT L POS NEG
.ENDS
***************************************
.SUBCKT aoi22 D0 S Y D1 GND VDD
** N=10 EP=6 IP=0 FDC=10
M0 9 D0 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.425e-13 AS=2.45e-13 PD=5.7e-07 PS=1.48e-06 $X=1380 $Y=-3795 $D=0
M1 Y 8 9 GND N_18 L=1.8e-07 W=5e-07 AD=1.2875e-13 AS=1.425e-13 PD=5.15e-07 PS=5.7e-07 $X=2130 $Y=-3795 $D=0
M2 10 D1 Y GND N_18 L=1.8e-07 W=5e-07 AD=1.3875e-13 AS=1.2875e-13 PD=5.55e-07 PS=5.15e-07 $X=2825 $Y=-3795 $D=0
M3 GND S 10 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.3875e-13 PD=5.1e-07 PS=5.55e-07 $X=3560 $Y=-3795 $D=0
M4 8 S GND GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=4250 $Y=-3795 $D=0
M5 5 D0 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=2.85e-13 AS=5.15e-13 PD=5.7e-07 PS=2.03e-06 $X=1380 $Y=-2130 $D=1
M6 Y S 5 VDD P_18 L=1.8e-07 W=1e-06 AD=2.575e-13 AS=2.85e-13 PD=5.15e-07 PS=5.7e-07 $X=2130 $Y=-2130 $D=1
M7 5 D1 Y VDD P_18 L=1.8e-07 W=1e-06 AD=2.775e-13 AS=2.575e-13 PD=5.55e-07 PS=5.15e-07 $X=2825 $Y=-2130 $D=1
M8 VDD 8 5 VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=2.775e-13 PD=5.1e-07 PS=5.55e-07 $X=3560 $Y=-2130 $D=1
M9 8 S VDD VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07 $X=4250 $Y=-2130 $D=1
.ENDS
***************************************
